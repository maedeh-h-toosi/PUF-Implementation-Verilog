`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:55:05 04/12/2021 
// Design Name: 
// Module Name:    RO 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RO1(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO2(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO3(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO4(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO5(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO6(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO7(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO8(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO9(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO10(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO11(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO12(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO13(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO14(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO15(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule

module RO16(input en,
			output out
    );

       (* S= "TRUE"*)(* ALLOW_COMBINATORIAL_LOOPS = "true", KEEP = "true" *) 
	    wire w1, w2, w3,w4,w5;  
		
		  
        and #1(w1, en, out);
        not #1(w2, w1);
        not #1(w3, w2);
        not #1(w4,w3);
        not #1(w5, w4);
        not #1(out, w5);
		  
endmodule